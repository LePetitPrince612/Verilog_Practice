module top_module(
    input               clk,
    input               x,
    output              z
    );

    
