module top_module(
    input               clk,
    input               L,
    input               r_in,
    input               q_in,
    output reg          Q
    );

    wire w;
    assign w = L? r_in : q_in;

    always_ff @(posedge clk) begin
        Q <= w;
    end

endmodule
